** sch_path: /home/Joerdson/LC_VCO.sch
**.subckt LC_VCO LON2 LOP2 VCC2 ICC2 GND VCTR2
*.iopin LON2
*.iopin LOP2
*.iopin VCC2
*.iopin ICC2
*.iopin VCTR2
*.iopin GND

XMN3 LOP2 LON2 net5 GND sg13_lv_nmos w=40.0u l=0.13u ng=5 m=1
XMN4 LON2 LOP2 net5 GND sg13_lv_nmos w=40.0u l=0.13u ng=5 m=1
XMN1 ICC2 ICC2 GND GND sg13_lv_nmos w=120.0u l=0.13u ng=15 m=1
XMN2 net5 ICC2 GND GND sg13_lv_nmos w=120.0u l=0.13u ng=15 m=1
XC1 VCC2 LOP2 cap_cmim w=8.73e-6 l=9.42e-6 m=1
XR1 LOP2 VCC2 rppd w=10.77e-6 l=8.92e-6 m=1 b=0
XC2 VCC2 LON2 cap_cmim w=8.73e-6 l=9.42e-6 m=1
XR2 LON2 VCC2 rppd w=10.77e-6 l=8.92e-6 m=1 b=0
L1 VCC2 LOP2 2.006n m=1
L2 VCC2 LON2 2.006n m=1
XCvar LOP2 VCTR2 LON2 net5 sg13_hv_svaricap W=9.74e-6 L=0.8e-6 Nx=2

**.ends
.end
